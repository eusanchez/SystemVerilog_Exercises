interface fizzbuzz_if (input logic clk);
    logic resetn;
    logic fizz;
    logic buzz;
    logic fizzbuzz;
endinterface //fizzbuzz_if 